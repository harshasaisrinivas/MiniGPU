`default_nettype none
`timescale 1ns/1ns
//Load-Store Unit
//Handles asynchronous memory load and store operations ans waits for response
//Each thread has its own LSU
//LDR, STR instructions are executed here
module lsu(
	input wire clk,
	input wire reset,
	input wire enable,
	//If current block has less threads than block size, some LSU will be inactive
	
	//State
	input reg[2:0] core_state,
	
	//Memory Control Signal
	input reg decoded_mem_read_enable,
	input reg decoded_mem_write_enable,
	
	//Registers
	input reg[7:0] rs,
	input reg[7:0] rt,
	
	//Data Memory
	output reg mem_read_valid,
	output reg[7:0] mem_read_address,
	input reg mem_read_ready,
	input reg[7:0] mem_read_data,
	output reg mem_write_valid,
	output reg[7:0] mem_write_address,
	output reg[7:0] mem_write_data,
	input reg mem_write_ready,
	
	//LSU outputs
	output reg[1:0] lsu_state,
	output reg[7:0] lsu_out
	);
	localparam IDLE = 2'b00, REQUESTING = 2'b01, WAITING = 2'b10, DONE = 2'b11;
	always@(posedge clk) begin
		if (reset) begin
			lsu_state <= IDLE;
			lsu_out <= 0;
			mem_read_valid <= 0;
			mem_read_address <= 0;
			mem_write_valid <= 0;
			mem_write_address <= 0;
			mem_write_data <=0;
			end
		else if(enable) begin
			//If memory read enable is triggered(LDR)
			if(decoded_mem_read_enable) begin
				case(lsu_state)
					IDLE: begin
					// Only read when core_state = REQUEST
						if(core_state == 3'b011) begin
							lsu_state <= REQUESTING;
						end
					end
					REQUESTING: begin
						mem_read_valid <= 1;
						mem_read_address <= rs;
						lsu_state <= WAITING;
					end
					WAITING: begin
						if(mem_read_ready == 1) begin
							mem_read_valid <= 0;
							lsu_out <= mem_read_data;
							lsu_state <= DONE;
						end
					end
					DONE: begin
						//Reset when core_state = UPDATE
						if(core_state == 3'b110) begin
							lsu_state <= IDLE;
						end
					end
				endcase
			end
			
			//If memory write enable is triggered(STR)
			if(decoded_mem_write_enable) begin
				case(lsu_state)
					IDLE: begin
						//Only write when core_state = REQUEST
						if(core_state == 3'b011) begin 
							lsu_state <= REQUESTING;
						end
					end
					REQUESTING: begin
						mem_write_valid <= 1;
						mem_write_address <= rs;
						mem_write_data <= rt;
						lsu_state <= WAITING;
					end
					WAITING: begin
						if(mem_write_ready) begin
							mem_write_valid <= 0;
							lsu_state <= DONE;
						end
					end
					DONE: begin
						//Reset when core_state = UPDATE
						if(core_state == 3'b1110) begin
							lsu_state <= IDLE;
						end
					end
				endcase
			end
		end
	end
endmodule
